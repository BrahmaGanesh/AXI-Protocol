package axi_pkg;

    `include "uvm_macros.svh"

    `include "axi_d"

endpackage