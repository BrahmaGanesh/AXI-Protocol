class axi_driver extends uvm_driver #(axi_transaction);
    `uvm_component_utils(axi_driver)

    virtual axi_interface vif;
    axi_transaction tr;

    function new(string name="axi_driver",uvm_component parent=null);
        super.new(name,parent);
    endfunction

    function void build_phase(uvm_phase phase);
        super.build_phase(phase);

        if(!uvm_config_db#(virtual axi_interface)::get(this,"","vif",vif))
            `uvm_fatal("DRV","axi_interface is not set")
    endfunction

    task run_phase(uvm_phase phase);
        forever begin
            seq_item_port.get_next_item(tr);
            if(tr.wr_en)begin
                vif.awvalid <= 1;
                vif.awaddr <= tr.awaddr;
                do @(posedge vif.clk);
                while(!vif.awready);
                vif.awvalid <= 0;

                vif.wdata <= tr.wdata;
                vif.wvalid <= 1;
                @(posedge vif.clk);
                wait(vif.wready);
                vif.wvalid <= 0;

                vif.bready <= 1;
                @(posedge vif.clk);
                wait(vif.bvalid);
                vif.bready <= 0;
                
                `uvm_info("DRV", $sformatf("Write transaction to address %0h with data %0h", tr.awaddr, tr.wdata), UVM_MEDIUM)
            end
            else begin
                vif.araddr <= tr.araddr;
                vif.arvalid <= 1;
                @(posedge vif.clk);
                wait(vif.arready);
                vif.arvalid <= 0;

                vif.rready <= 1;
                @(posedge vif.clk);
                wait(vif.rvalid);
                vif.rready <= 0;

                `uvm_info("DRV", $sformatf("Read transaction from address %0h", tr.araddr), UVM_MEDIUM)
            end
            seq_item_port.item_done();
            #1;
        end
    endtask
endclass
